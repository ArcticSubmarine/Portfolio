library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
library AESLibrary;
use AESLibrary.state_definition_package.all;


entity InvAESRound is 
	port (	clock_i			: in std_logic;	--Signal d'horloge
		currentKey_i		: in bit128;	--Clé courrante
		currentText_i		: in bit128;	--Texte courrant
		enableInvMixColumns_i	: in std_logic;	--Signal autorisant InvMixColumns
		enableRoundComputing_i	: in std_logic;	--Signal autorisant RoundComputing
		resetb_i		: in std_logic;	--Signal de reset
		data_o			: out bit128);	--Sortie
end entity;


architecture InvAESRound_arch of InvAESRound is
	component AddRoundKey is
		port (	AddRoundKey_i 	: in type_state;	--Clé courrante
			Expansion_key_i : in type_state;	--Texte courrant
			AddRoundKey_o 	: out type_state);
	end component AddRoundKey;

	component InvShiftRows is
	port (	InvShiftRows_i : in type_state;
		InvShiftRows_o : out type_state);
	end component InvShiftRows;

	component InvSubBytes is 
	port (	InvSubBytes_i : in type_state;
		InvSubBytes_o : out type_state);
	end component InvSubBytes;

	component InvMixColumns is
		port (	InvMixColumns_i : in type_state;
			InvMixColumns_o : out type_state);
	end component InvMixColumns;

	type state is (initialisation, debut, boucle, fin);	
	signal etat_actuel, etat_futur : state;	--Etat d'avancement de l'algorithme

	signal currentKey_s		: type_state;
	signal currentText_s		: type_state;
	signal AddRoundKey_i_s		: type_state;
	signal Expansion_key_i_s	: type_state;
	signal AddRoundKey_o_s		: type_state;
	signal InvShiftRows_i_s		: type_state;
	signal InvShiftRows_o_s		: type_state;
	signal InvSubBytes_i_s		: type_state;
	signal InvSubBytes_o_s		: type_state;
	signal InvMixColumns_i_s	: type_state;
	signal InvMixColumns_o_s	: type_state;


	begin
		DUT : AddRoundKey
		port map (	AddRoundKey_i 		=> AddRoundKey_i_s,	--Clé courrante
				Expansion_key_i 	=> Expansion_key_i_s,	--Texte courrant
				AddRoundKey_o 		=> AddRoundKey_o_s);

		DUT1 : InvSubBytes
		port map (	InvSubBytes_i	=> InvSubBytes_i_s,
				InvSubBytes_o	=> InvSubBytes_o_s);

		DUT2 : InvShiftRows
		port map (	InvShiftRows_i	=> InvShiftRows_i_s,
				InvShiftRows_o	=> InvShiftRows_o_s);

		DUT3 : InvMixColumns
		port map (	InvMixColumns_i	=> InvMixColumns_i_s,
				InvMixColumns_o	=> InvMixColumns_o_s);

	
		P0 : process (clock_i, resetb_i)	--Cas reset
		begin
			if resetb_i = '1' then etat_actuel <= initialisation;
			elsif clock_i'event and clock_i = '1' then 
				etat_actuel <= etat_futur;
			end if;
		end process P0;


		P1 : process (etat_actuel, enableInvMixColumns_i, enableRoundComputing_i)
		begin
			case etat_actuel is
				when initialisation =>
					if enableRoundComputing_i = '1' then etat_futur <= debut;
					else 
						etat_futur <= initialisation;
					end if;
	
				when debut => 
					if enableInvMixColumns_i = '1' then
						etat_futur <= boucle;
					else 
				  		etat_futur <= debut;
					end if;
	
				when boucle => 
					if enableRoundComputing_i = '0' then 
					 	etat_futur <= fin;
					else 
					   	etat_futur <= boucle;
					end if;
		
				when fin =>
					if resetb_i = '0' then
					 	etat_futur <= fin;
					else 
					  	etat_futur <= initialisation;
					end if;
			end case;
		end process P1;
		
		P2 : process (etat_actuel)
		begin 
			case etat_actuel is 
				when initialisation =>
					currentText_s(0)(0) <= currentText_i(7	downto 0);
					currentText_s(0)(1) <= currentText_i(15 downto 8);
					currentText_s(0)(2) <= currentText_i(23 downto 16);
					currentText_s(0)(3) <= currentText_i(31 downto 24);
					currentText_s(1)(0) <= currentText_i(39 downto 32);
					currentText_s(1)(1) <= currentText_i(47 downto 40);
					currentText_s(1)(2) <= currentText_i(55 downto 48);
					currentText_s(1)(3) <= currentText_i(63 downto 56);
					currentText_s(2)(0) <= currentText_i(71 downto 64);
					currentText_s(2)(1) <= currentText_i(79 downto 72);
					currentText_s(2)(2) <= currentText_i(87 downto 80);
					currentText_s(2)(3) <= currentText_i(95 downto 88);
					currentText_s(3)(0) <= currentText_i(103 downto 96);
					currentText_s(3)(1) <= currentText_i(111 downto 104);
					currentText_s(3)(2) <= currentText_i(119 downto 112);
					currentText_s(3)(3) <= currentText_i(127 downto 120);

					currentKey_s(0)(0) <= currentKey_i(7 downto 0);
					currentKey_s(0)(1) <= currentKey_i(15 downto 8);
					currentKey_s(0)(2) <= currentKey_i(23 downto 16);
					currentKey_s(0)(3) <= currentKey_i(31 downto 24);
					currentKey_s(1)(0) <= currentKey_i(39 downto 32);
					currentKey_s(1)(1) <= currentKey_i(47 downto 40);
					currentKey_s(1)(2) <= currentKey_i(55 downto 48);
					currentKey_s(1)(3) <= currentKey_i(63 downto 56);
					currentKey_s(2)(0) <= currentKey_i(71 downto 64);
					currentKey_s(2)(1) <= currentKey_i(79 downto 72);
					currentKey_s(2)(2) <= currentKey_i(87 downto 80);
					currentKey_s(2)(3) <= currentKey_i(95 downto 88);
					currentKey_s(3)(0) <= currentKey_i(103 downto 96);
					currentKey_s(3)(1) <= currentKey_i(111 downto 104);
					currentKey_s(3)(2) <= currentKey_i(119 downto 112);
					currentKey_s(3)(3) <= currentKey_i(127 downto 120);
			
				when debut =>
					AddRoundKey_i_s 	<= currentText_s;
					Expansion_key_i_s	<= currentKey_s;

				when boucle =>
					InvSubBytes_i_s		<= AddRoundKey_o_s;
					InvShiftRows_i_s	<= InvSubBytes_o_s;
					InvMixColumns_i_s	<= InvShiftRows_o_s;
					AddRoundKey_i_s		<= InvMixColumns_o_s;
				
				when fin =>		
					InvSubBytes_i_s		<= AddRoundKey_o_s;
					InvShiftRows_i_s	<= InvSubBytes_o_s;
					AddRoundKey_i_s		<= InvShiftRows_o_s;

					data_o(7 downto 0)	<= AddRoundKey_o_s(0)(0);
					data_o(15 downto 8)	<= AddRoundKey_o_s(0)(1);
					data_o(23 downto 16)	<= AddRoundKey_o_s(0)(2);
					data_o(31 downto 24)	<= AddRoundKey_o_s(0)(3);		
					data_o(39 downto 32)	<= AddRoundKey_o_s(1)(0);
					data_o(47 downto 40)	<= AddRoundKey_o_s(1)(1);
					data_o(55 downto 48)	<= AddRoundKey_o_s(1)(2);
					data_o(63 downto 56)	<= AddRoundKey_o_s(1)(3);
					data_o(71 downto 64)	<= AddRoundKey_o_s(2)(0);
					data_o(79 downto 72)	<= AddRoundKey_o_s(2)(1);
					data_o(87 downto 80)	<= AddRoundKey_o_s(2)(2);
					data_o(95 downto 88)	<= AddRoundKey_o_s(2)(3);
					data_o(103 downto 96)	<= AddRoundKey_o_s(3)(0);
					data_o(111 downto 104)	<= AddRoundKey_o_s(3)(1);
					data_o(119 downto 112)	<= AddRoundKey_o_s(3)(2);
					data_o(127 downto 120)	<= AddRoundKey_o_s(3)(3);
					
			end case;	
		end process P2;

end architecture;
